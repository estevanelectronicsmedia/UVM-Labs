// Activity 01:

`include "uvm_macros.svh"
import uvm_pkg::*;
 
module tb;
  initial begin
    `uvm_info("Testbench", $sformatf("First RTL Code : %0s","Half Adder"), UVM_NONE);
  end
  
endmodule
